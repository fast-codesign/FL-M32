/*
 *  Project:            timelyRV_v0.1 -- a RISCV-32I SoC.
 *  Module name:        timelyRV_core, i.e., a simplified picorv32.
 *  Description:        RISCV-32I core.
 *  Last updated date:  2022.04.02.
 *
 *  Copyright (C) 2021-2022 Junnan Li <lijunnan@nudt.edu.cn>.
 *  Copyright and related rights are licensed under the MIT license.
 *
 */

`timescale 1 ns / 1 ps

/***************************************************************
 * picorv32
 ***************************************************************/

module picorv32_simplified #(
  parameter [ 0:0] ENABLE_COUNTERS = 1,
  parameter [ 0:0] ENABLE_COUNTERS64 = 1,
  parameter [ 0:0] ENABLE_REGS_16_31 = 1,
  parameter [ 0:0] ENABLE_REGS_DUALPORT = 1,
  parameter [ 0:0] LATCHED_MEM_RDATA = 0,
  parameter [ 0:0] TWO_STAGE_SHIFT = 1,
  parameter [ 0:0] BARREL_SHIFTER = 0,
  parameter [ 0:0] TWO_CYCLE_COMPARE = 0,
  parameter [ 0:0] TWO_CYCLE_ALU = 0,
  parameter [ 0:0] COMPRESSED_ISA = 0,
  parameter [ 0:0] CATCH_MISALIGN = 1,
  parameter [ 0:0] CATCH_ILLINSN = 1,
  parameter [ 0:0] ENABLE_PCPI = 0,
  parameter [ 0:0] ENABLE_MUL = 0,
  parameter [ 0:0] ENABLE_FAST_MUL = 0,
  parameter [ 0:0] ENABLE_DIV = 0,
  parameter [ 0:0] ENABLE_IRQ = 1,
  parameter [ 0:0] ENABLE_IRQ_QREGS = 1,
  parameter [ 0:0] ENABLE_IRQ_TIMER = 1,
  parameter [ 0:0] ENABLE_TRACE = 0,
  parameter [ 0:0] REGS_INIT_ZERO = 0,
  parameter [31:0] MASKED_IRQ = 32'h 0000_0000,
  parameter [31:0] LATCHED_IRQ = 32'h ffff_ffff,
  parameter [31:0] PROGADDR_RESET = 32'h 0000_0000,
  parameter [31:0] PROGADDR_IRQ = 32'h 0000_0010,
  parameter [31:0] STACKADDR = 32'h ffff_ffff
) (
  input clk, resetn,
  output reg trap,

  output reg        mem_valid,
  output reg        mem_instr,
  input             mem_ready,

  output reg [31:0] mem_addr,
  output reg [31:0] mem_wdata,
  output reg [ 3:0] mem_wstrb,
  input      [31:0] mem_rdata,

  // Look-Ahead Interface
  output            mem_la_read,
  output            mem_la_write,
  output     [31:0] mem_la_addr,
  output reg [31:0] mem_la_wdata,
  output reg [ 3:0] mem_la_wstrb,

  // IRQ Interface
  input      [31:0] irq,
  output reg [31:0] eoi,

  // Trace Interface
  output reg        trace_valid,
  output reg [35:0] trace_data
);
  localparam integer irq_timer = 0;
  localparam integer irq_ebreak = 1;
  localparam integer irq_buserror = 2;

  localparam integer irqregs_offset = ENABLE_REGS_16_31 ? 32 : 16;
  localparam integer regfile_size = (ENABLE_REGS_16_31 ? 32 : 16) + 4*ENABLE_IRQ*ENABLE_IRQ_QREGS;
  localparam integer regindex_bits = (ENABLE_REGS_16_31 ? 5 : 4) + ENABLE_IRQ*ENABLE_IRQ_QREGS;


  localparam [35:0] TRACE_BRANCH = {4'b 0001, 32'b 0};
  localparam [35:0] TRACE_ADDR   = {4'b 0010, 32'b 0};
  localparam [35:0] TRACE_IRQ    = {4'b 1000, 32'b 0};

  // for cpu irq disable
  localparam [31:0] SYS_MASKED_IRQ = 32'h ffff_fff9;

  reg [63:0] count_cycle, count_instr;
  
  //* reg_pc used for jal, jalr, branch instructions;
  //* reg_next_pc for reading instruction as address;
  //* reg_op1 is the first operation register;
  //* reg_op2 is the second operation register;
  //* reg_out is the result of not alu instructions, e.g., jalr, branch;
  //* reg_sh for shift;
  reg [31:0] reg_pc, reg_next_pc, reg_op1, reg_op2, reg_out;
  reg [4:0] reg_sh;

  //* next_pc used as address to read instruction;
  wire [31:0] next_pc;

  reg irq_delay;
  reg irq_active;
  reg [31:0] irq_mask;
  reg irq_on;
  reg [31:0] irq_pending;
  reg [31:0] timer, timer_conf;

  //* cpu regs;
  reg [31:0] cpuregs [0:regfile_size-1];
  integer i;
  initial begin
    if (REGS_INIT_ZERO) begin
      for (i = 0; i < regfile_size; i = i+1)
        cpuregs[i] = 0;
    end
  end

  //* Memory Interface
  reg [1:0] mem_state;    //* state of reading/writing memory;
  reg [1:0] mem_wordsize;   //* number of bytes to read/write;
  reg [31:0] mem_rdata_word;  //* rdata of data;
  reg [31:0] mem_rdata_q;   //* store mem_rdata for decoding at the second stage;
  reg mem_do_prefetch;    //* to prefetch instruction;
  reg mem_do_rinst;     //* to read instruction;
  reg mem_do_rdata;     //* to read data;
  reg mem_do_wdata;     //* to write data;

  
  //* mem_rdata is valid;
  wire mem_xfer;
  assign mem_xfer = mem_valid && mem_ready;

  //* finish memory reading/writing (include prefetch has received mem_do_rinst);
  wire mem_done = resetn && ((mem_xfer && |mem_state && (mem_do_rinst || mem_do_rdata || mem_do_wdata)) || (&mem_state && mem_do_rinst));

  //* mem_la_write/read/addr is valid when mem_do_wdata/rinst/prefetch/rdata is valid;
  assign mem_la_write = resetn && !mem_state && mem_do_wdata;
  assign mem_la_read = resetn && (!mem_state && (mem_do_rinst || mem_do_prefetch || mem_do_rdata));
  assign mem_la_addr = (mem_do_prefetch || mem_do_rinst) ? {next_pc[31:2], 2'b00} : {reg_op1[31:2], 2'b00};
  
  //* used for first-stage decode, = mem_rdata (for rinst) or = mem_rdata_q (for instr_prefetch)
  wire [31:0] mem_rdata_latched;
  assign mem_rdata_latched = (mem_xfer || LATCHED_MEM_RDATA) ? mem_rdata : mem_rdata_q;

  //* write/read according to mem_wordsize
  always @* begin
    (* full_case *)
    case (mem_wordsize)
      0: begin
        mem_la_wdata = reg_op2;
        mem_la_wstrb = 4'b1111;
        mem_rdata_word = mem_rdata;
      end
      1: begin
        mem_la_wdata = {2{reg_op2[15:0]}};
        mem_la_wstrb = reg_op1[1] ? 4'b1100 : 4'b0011;
        case (reg_op1[1])
          1'b0: mem_rdata_word = {16'b0, mem_rdata[15: 0]};
          1'b1: mem_rdata_word = {16'b0, mem_rdata[31:16]};
        endcase
      end
      2: begin
        mem_la_wdata = {4{reg_op2[7:0]}};
        mem_la_wstrb = 4'b0001 << reg_op1[1:0];
        case (reg_op1[1:0])
          2'b00: mem_rdata_word = {24'b0, mem_rdata[ 7: 0]};
          2'b01: mem_rdata_word = {24'b0, mem_rdata[15: 8]};
          2'b10: mem_rdata_word = {24'b0, mem_rdata[23:16]};
          2'b11: mem_rdata_word = {24'b0, mem_rdata[31:24]};
        endcase
      end
    endcase
  end

  always @(posedge clk) begin
    if (mem_xfer) begin
      mem_rdata_q <= mem_rdata;
    end
  end

  //* assign memory interface signals;
  always @(posedge clk) begin
    if (!resetn || trap) begin
      if (!resetn)
        mem_state <= 0;
      if (!resetn || mem_ready)
        mem_valid <= 0;
    end else begin
      if (mem_la_read || mem_la_write) begin
        mem_addr <= mem_la_addr;
        mem_wstrb <= mem_la_wstrb & {4{mem_la_write}};
      end
      if (mem_la_write) begin
        mem_wdata <= mem_la_wdata;
      end
      case (mem_state)
        0: begin
          if (mem_do_prefetch || mem_do_rinst || mem_do_rdata) begin
            mem_valid <= 1;
            mem_instr <= mem_do_prefetch || mem_do_rinst;
            mem_wstrb <= 0;
            mem_state <= 1;
          end
          if (mem_do_wdata) begin
            mem_valid <= 1;
            mem_instr <= 0;
            mem_state <= 2;
          end
        end
        1: begin
          if (mem_xfer) begin
            mem_valid <= 0;
            mem_state <= mem_do_rinst || mem_do_rdata ? 0 : 3;
          end
        end
        2: begin
          if (mem_xfer) begin
            mem_valid <= 0;
            mem_state <= 0;
          end
        end
        3: begin
          if (mem_do_rinst) begin
            mem_state <= 0;
          end
        end
      endcase
    end

  end


  // Instruction Decoder

  reg instr_lui, instr_auipc, instr_jal, instr_jalr;
  reg instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu;
  reg instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw;
  reg instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai;
  reg instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and;
  reg instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh, instr_ecall_ebreak;
  reg instr_getq, instr_setq, instr_retirq, instr_maskirq, instr_waitirq, instr_timer, instr_ctlirq;
  wire instr_trap;

  reg [regindex_bits-1:0] decoded_rd, decoded_rs1, decoded_rs2;
  reg [31:0] decoded_imm, decoded_imm_j;
  reg decoder_trigger;
  reg decoder_trigger_q;
  reg decoder_pseudo_trigger;
  reg decoder_pseudo_trigger_q;
  // reg compressed_instr;

  reg is_lui_auipc_jal;
  reg is_lb_lh_lw_lbu_lhu;
  reg is_slli_srli_srai;
  reg is_jalr_addi_slti_sltiu_xori_ori_andi;
  reg is_sb_sh_sw;
  reg is_sll_srl_sra;
  reg is_lui_auipc_jal_jalr_addi_add_sub;
  reg is_slti_blt_slt;
  reg is_sltiu_bltu_sltu;
  reg is_beq_bne_blt_bge_bltu_bgeu;
  reg is_lbu_lhu_lw;
  reg is_alu_reg_imm;
  reg is_alu_reg_reg;
  reg is_compare;

  assign instr_trap = CATCH_ILLINSN && !{instr_lui, instr_auipc, instr_jal, instr_jalr,
      instr_beq, instr_bne, instr_blt, instr_bge, instr_bltu, instr_bgeu,
      instr_lb, instr_lh, instr_lw, instr_lbu, instr_lhu, instr_sb, instr_sh, instr_sw,
      instr_addi, instr_slti, instr_sltiu, instr_xori, instr_ori, instr_andi, instr_slli, instr_srli, instr_srai,
      instr_add, instr_sub, instr_sll, instr_slt, instr_sltu, instr_xor, instr_srl, instr_sra, instr_or, instr_and,
      instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh,
      instr_getq, instr_setq, instr_retirq, instr_maskirq, instr_waitirq, instr_timer, instr_ctlirq};

  wire is_rdcycle_rdcycleh_rdinstr_rdinstrh;
  assign is_rdcycle_rdcycleh_rdinstr_rdinstrh = |{instr_rdcycle, instr_rdcycleh, instr_rdinstr, instr_rdinstrh};

  //* two-stage decode;
  always @(posedge clk) begin
    //* second stage;
    is_lui_auipc_jal <= |{instr_lui, instr_auipc, instr_jal};
    is_lui_auipc_jal_jalr_addi_add_sub <= |{instr_lui, instr_auipc, instr_jal, instr_jalr, instr_addi, instr_add, instr_sub};
    is_slti_blt_slt <= |{instr_slti, instr_blt, instr_slt};
    is_sltiu_bltu_sltu <= |{instr_sltiu, instr_bltu, instr_sltu};
    is_lbu_lhu_lw <= |{instr_lbu, instr_lhu, instr_lw};
    is_compare <= |{is_beq_bne_blt_bge_bltu_bgeu, instr_slti, instr_slt, instr_sltiu, instr_sltu};

    //* first stage;
    if (mem_do_rinst && mem_done) begin
      instr_lui     <= mem_rdata_latched[6:0] == 7'b0110111;
      instr_auipc   <= mem_rdata_latched[6:0] == 7'b0010111;
      instr_jal     <= mem_rdata_latched[6:0] == 7'b1101111;
      instr_jalr    <= mem_rdata_latched[6:0] == 7'b1100111 && mem_rdata_latched[14:12] == 3'b000;
      instr_retirq  <= mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000010 && ENABLE_IRQ;
      instr_waitirq <= mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000100 && ENABLE_IRQ;

      is_beq_bne_blt_bge_bltu_bgeu <= mem_rdata_latched[6:0] == 7'b1100011;
      is_lb_lh_lw_lbu_lhu          <= mem_rdata_latched[6:0] == 7'b0000011;
      is_sb_sh_sw                  <= mem_rdata_latched[6:0] == 7'b0100011;
      is_alu_reg_imm               <= mem_rdata_latched[6:0] == 7'b0010011;
      is_alu_reg_reg               <= mem_rdata_latched[6:0] == 7'b0110011;

      { decoded_imm_j[31:20], decoded_imm_j[10:1], decoded_imm_j[11], decoded_imm_j[19:12], decoded_imm_j[0] } <= $signed({mem_rdata_latched[31:12], 1'b0});

      decoded_rd <= mem_rdata_latched[11:7];
      decoded_rs1 <= mem_rdata_latched[19:15];
      decoded_rs2 <= mem_rdata_latched[24:20];

      if (mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000000 && ENABLE_IRQ && ENABLE_IRQ_QREGS)
        decoded_rs1[regindex_bits-1] <= 1; // instr_getq

      if (mem_rdata_latched[6:0] == 7'b0001011 && mem_rdata_latched[31:25] == 7'b0000010 && ENABLE_IRQ)
        decoded_rs1 <= ENABLE_IRQ_QREGS ? irqregs_offset : 3; // instr_retirq

      // compressed_instr <= 0;
    end

    //* second stage;
    if (decoder_trigger && !decoder_pseudo_trigger) begin

      instr_beq   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b000;
      instr_bne   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b001;
      instr_blt   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b100;
      instr_bge   <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b101;
      instr_bltu  <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b110;
      instr_bgeu  <= is_beq_bne_blt_bge_bltu_bgeu && mem_rdata_q[14:12] == 3'b111;

      instr_lb    <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b000;
      instr_lh    <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b001;
      instr_lw    <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b010;
      instr_lbu   <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b100;
      instr_lhu   <= is_lb_lh_lw_lbu_lhu && mem_rdata_q[14:12] == 3'b101;

      instr_sb    <= is_sb_sh_sw && mem_rdata_q[14:12] == 3'b000;
      instr_sh    <= is_sb_sh_sw && mem_rdata_q[14:12] == 3'b001;
      instr_sw    <= is_sb_sh_sw && mem_rdata_q[14:12] == 3'b010;

      instr_addi  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b000;
      instr_slti  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b010;
      instr_sltiu <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b011;
      instr_xori  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b100;
      instr_ori   <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b110;
      instr_andi  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b111;

      instr_slli  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000;
      instr_srli  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000;
      instr_srai  <= is_alu_reg_imm && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000;

      instr_add   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b000 && mem_rdata_q[31:25] == 7'b0000000;
      instr_sub   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b000 && mem_rdata_q[31:25] == 7'b0100000;
      instr_sll   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000;
      instr_slt   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b010 && mem_rdata_q[31:25] == 7'b0000000;
      instr_sltu  <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b011 && mem_rdata_q[31:25] == 7'b0000000;
      instr_xor   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b100 && mem_rdata_q[31:25] == 7'b0000000;
      instr_srl   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000;
      instr_sra   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000;
      instr_or    <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b110 && mem_rdata_q[31:25] == 7'b0000000;
      instr_and   <= is_alu_reg_reg && mem_rdata_q[14:12] == 3'b111 && mem_rdata_q[31:25] == 7'b0000000;

      instr_rdcycle  <= ((mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11000000000000000010) ||
                         (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11000000000100000010)) && ENABLE_COUNTERS;
      instr_rdcycleh <= ((mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11001000000000000010) ||
                         (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11001000000100000010)) && ENABLE_COUNTERS && ENABLE_COUNTERS64;
      instr_rdinstr  <=  (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11000000001000000010) && ENABLE_COUNTERS;
      instr_rdinstrh <=  (mem_rdata_q[6:0] == 7'b1110011 && mem_rdata_q[31:12] == 'b11001000001000000010) && ENABLE_COUNTERS && ENABLE_COUNTERS64;

      instr_ecall_ebreak <= (mem_rdata_q[6:0] == 7'b1110011 && !mem_rdata_q[31:21] && !mem_rdata_q[19:7]);

      instr_getq    <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000000 && ENABLE_IRQ && ENABLE_IRQ_QREGS;
      instr_setq    <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000001 && ENABLE_IRQ && ENABLE_IRQ_QREGS;
      instr_maskirq <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000011 && ENABLE_IRQ;
      instr_timer   <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000101 && ENABLE_IRQ && ENABLE_IRQ_TIMER;
      instr_ctlirq  <= mem_rdata_q[6:0] == 7'b0001011 && mem_rdata_q[31:25] == 7'b0000110 && ENABLE_IRQ;

      is_slli_srli_srai <= is_alu_reg_imm && |{
        mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000,
        mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000,
        mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000
      };

      is_jalr_addi_slti_sltiu_xori_ori_andi <= instr_jalr || is_alu_reg_imm && |{
        mem_rdata_q[14:12] == 3'b000,
        mem_rdata_q[14:12] == 3'b010,
        mem_rdata_q[14:12] == 3'b011,
        mem_rdata_q[14:12] == 3'b100,
        mem_rdata_q[14:12] == 3'b110,
        mem_rdata_q[14:12] == 3'b111
      };

      is_sll_srl_sra <= is_alu_reg_reg && |{
        mem_rdata_q[14:12] == 3'b001 && mem_rdata_q[31:25] == 7'b0000000,
        mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0000000,
        mem_rdata_q[14:12] == 3'b101 && mem_rdata_q[31:25] == 7'b0100000
      };

      is_lui_auipc_jal_jalr_addi_add_sub <= 0;
      is_compare <= 0;

      (* parallel_case *)
      case (1'b1)
        instr_jal:
          decoded_imm <= decoded_imm_j;
        |{instr_lui, instr_auipc}:
          decoded_imm <= mem_rdata_q[31:12] << 12;
        |{instr_jalr, is_lb_lh_lw_lbu_lhu, is_alu_reg_imm}:
          decoded_imm <= $signed(mem_rdata_q[31:20]);
        is_beq_bne_blt_bge_bltu_bgeu:
          decoded_imm <= $signed({mem_rdata_q[31], mem_rdata_q[7], mem_rdata_q[30:25], mem_rdata_q[11:8], 1'b0});
        is_sb_sh_sw:
          decoded_imm <= $signed({mem_rdata_q[31:25], mem_rdata_q[11:7]});
        default:
          decoded_imm <= 1'bx;
      endcase
    end

    if (!resetn) begin
      is_beq_bne_blt_bge_bltu_bgeu <= 0;
      is_compare <= 0;

      instr_beq   <= 0;
      instr_bne   <= 0;
      instr_blt   <= 0;
      instr_bge   <= 0;
      instr_bltu  <= 0;
      instr_bgeu  <= 0;

      instr_addi  <= 0;
      instr_slti  <= 0;
      instr_sltiu <= 0;
      instr_xori  <= 0;
      instr_ori   <= 0;
      instr_andi  <= 0;

      instr_add   <= 0;
      instr_sub   <= 0;
      instr_sll   <= 0;
      instr_slt   <= 0;
      instr_sltu  <= 0;
      instr_xor   <= 0;
      instr_srl   <= 0;
      instr_sra   <= 0;
      instr_or    <= 0;
      instr_and   <= 0;
    end
  end


  // Main State Machine

  localparam cpu_state_trap   = 8'b10000000;
  localparam cpu_state_fetch  = 8'b01000000;
  localparam cpu_state_ld_rs1 = 8'b00100000;
  localparam cpu_state_ld_rs2 = 8'b00010000;
  localparam cpu_state_exec   = 8'b00001000;
  localparam cpu_state_shift  = 8'b00000100;
  localparam cpu_state_stmem  = 8'b00000010;
  localparam cpu_state_ldmem  = 8'b00000001;

  reg [7:0] cpu_state;
  reg [1:0] irq_state;  //* ?


  reg set_mem_do_rinst; //* to set mem_do_rinst;
  reg set_mem_do_rdata; //* to set mem_do_rdata;
  reg set_mem_do_wdata; //* to set mem_do_wdata;

  reg latched_store;    //* to write register( is '0' while branch miss 
              //*   jal instr or store instr);
  reg latched_stalu;    //* not branch, jal instruction;
  reg latched_branch;   //* branch (hit), jalr, jal;
  // reg latched_compr;
  reg latched_trace;
  reg latched_is_lu;    //* used at cpu_state_ldmem
  reg latched_is_lh;
  reg latched_is_lb;
  reg [regindex_bits-1:0] latched_rd; //* which register to wirte;

  reg [31:0] current_pc;  //* used to calculate reg_next_pc;
  assign next_pc = latched_store && latched_branch ? reg_out & ~1 : reg_next_pc;


  reg [31:0] next_irq_pending;
  reg do_waitirq;

  reg [31:0] alu_out, alu_out_q;  //* result of alu;
  reg alu_out_0, alu_out_0_q;   //* result of cmp;
  reg alu_wait, alu_wait_2;   //* usedw at cpu_stage_exec;

  reg [31:0] alu_add_sub;
  reg [31:0] alu_shl, alu_shr;
  reg alu_eq, alu_ltu, alu_lts;

  generate if (TWO_CYCLE_ALU) begin
    always @(posedge clk) begin
      alu_add_sub <= instr_sub ? reg_op1 - reg_op2 : reg_op1 + reg_op2;
      alu_eq <= reg_op1 == reg_op2;
      alu_lts <= $signed(reg_op1) < $signed(reg_op2);
      alu_ltu <= reg_op1 < reg_op2;
      alu_shl <= reg_op1 << reg_op2[4:0];
      alu_shr <= $signed({instr_sra || instr_srai ? reg_op1[31] : 1'b0, reg_op1}) >>> reg_op2[4:0];
    end
  end else begin
    always @* begin
      alu_add_sub = instr_sub ? reg_op1 - reg_op2 : reg_op1 + reg_op2;
      alu_eq = reg_op1 == reg_op2;
      alu_lts = $signed(reg_op1) < $signed(reg_op2);
      alu_ltu = reg_op1 < reg_op2;
      alu_shl = reg_op1 << reg_op2[4:0];
      alu_shr = $signed({instr_sra || instr_srai ? reg_op1[31] : 1'b0, reg_op1}) >>> reg_op2[4:0];
    end
  end endgenerate

  always @* begin
    alu_out_0 = 'bx;
    (* parallel_case, full_case *)
    case (1'b1)
      instr_beq:
        alu_out_0 = alu_eq;
      instr_bne:
        alu_out_0 = !alu_eq;
      instr_bge:
        alu_out_0 = !alu_lts;
      instr_bgeu:
        alu_out_0 = !alu_ltu;
      is_slti_blt_slt && (!TWO_CYCLE_COMPARE || !{instr_beq,instr_bne,instr_bge,instr_bgeu}):
        alu_out_0 = alu_lts;
      is_sltiu_bltu_sltu && (!TWO_CYCLE_COMPARE || !{instr_beq,instr_bne,instr_bge,instr_bgeu}):
        alu_out_0 = alu_ltu;
    endcase

    alu_out = 'bx;
    (* parallel_case, full_case *)
    case (1'b1)
      is_lui_auipc_jal_jalr_addi_add_sub:
        alu_out = alu_add_sub;
      is_compare:
        alu_out = alu_out_0;
      instr_xori || instr_xor:
        alu_out = reg_op1 ^ reg_op2;
      instr_ori || instr_or:
        alu_out = reg_op1 | reg_op2;
      instr_andi || instr_and:
        alu_out = reg_op1 & reg_op2;
      BARREL_SHIFTER && (instr_sll || instr_slli):
        alu_out = alu_shl;
      BARREL_SHIFTER && (instr_srl || instr_srli || instr_sra || instr_srai):
        alu_out = alu_shr;
    endcase
  end


  reg cpuregs_write;
  reg [31:0] cpuregs_wrdata;
  reg [31:0] cpuregs_rs1;
  reg [31:0] cpuregs_rs2;

  always @* begin
    cpuregs_write = 0;
    cpuregs_wrdata = 'bx;

    if (cpu_state == cpu_state_fetch) begin
      (* parallel_case *)
      case (1'b1)
        latched_branch: begin   // exclude branch／retirq instr, as latched_rd = 0;
          cpuregs_wrdata = reg_pc + 4;
          cpuregs_write = 1;
        end
        latched_store && !latched_branch: begin
          cpuregs_wrdata = latched_stalu ? alu_out_q : reg_out;
          cpuregs_write = 1;
        end
        ENABLE_IRQ && irq_state[0]: begin
          cpuregs_wrdata = reg_next_pc;
          cpuregs_write = 1;
        end
        ENABLE_IRQ && irq_state[1]: begin
          cpuregs_wrdata = irq_pending & ~irq_mask;
          cpuregs_write = 1;
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if (resetn && cpuregs_write && latched_rd)
      cpuregs[latched_rd] <= cpuregs_wrdata;
  end

  always @* begin
    cpuregs_rs1 = decoded_rs1 ? cpuregs[decoded_rs1] : 0;
    cpuregs_rs2 = decoded_rs2 ? cpuregs[decoded_rs2] : 0;
  end

  
  always @(posedge clk) begin
    trap <= 0;
    reg_sh <= 'bx;
    reg_out <= 'bx;
    set_mem_do_rinst = 0;
    set_mem_do_rdata = 0;
    set_mem_do_wdata = 0;

    alu_out_0_q <= alu_out_0;
    alu_out_q <= alu_out;

    alu_wait <= 0;
    alu_wait_2 <= 0;


    if (ENABLE_COUNTERS) begin
      count_cycle <= resetn ? count_cycle + 1 : 0;
      if (!ENABLE_COUNTERS64) count_cycle[63:32] <= 0;
    end else begin
      count_cycle <= 'bx;
      count_instr <= 'bx;
    end

    next_irq_pending = ENABLE_IRQ ? irq_pending & LATCHED_IRQ : 'bx;

    if (ENABLE_IRQ && ENABLE_IRQ_TIMER && timer) begin
      timer <= timer - 1;
      if (timer - 1 == 0) begin
        next_irq_pending[irq_timer] = 1;
        timer   <= timer_conf;
      end
    end

    if (ENABLE_IRQ) begin
      next_irq_pending = next_irq_pending | irq;
    end

    decoder_trigger <= mem_do_rinst && mem_done;
    decoder_trigger_q <= decoder_trigger;
    decoder_pseudo_trigger <= 0;
    decoder_pseudo_trigger_q <= decoder_pseudo_trigger;
    do_waitirq <= 0;

    trace_valid <= 0;

    if (!ENABLE_TRACE)
      trace_data <= 'bx;

    if (!resetn) begin
      reg_pc <= PROGADDR_RESET;
      reg_next_pc <= PROGADDR_RESET;
      if (ENABLE_COUNTERS)
        count_instr <= 0;
      latched_store <= 0;
      latched_stalu <= 0;
      latched_branch <= 0;
      latched_trace <= 0;
      latched_is_lu <= 0;
      latched_is_lh <= 0;
      latched_is_lb <= 0;
      irq_active <= 0;
      irq_delay <= 0;
      irq_mask <= ~0;
      irq_on <= 0;
      next_irq_pending = 0;
      irq_state <= 0;
      eoi <= 0;
      timer <= 0;
      timer_conf <= 0;
      if (~STACKADDR) begin
        latched_store <= 1;
        latched_rd <= 2;
        reg_out <= STACKADDR;
      end
      cpu_state <= cpu_state_fetch;
    end else
    (* parallel_case, full_case *)
    case (cpu_state)
      cpu_state_trap: begin
        trap <= 1;
      end

      cpu_state_fetch: begin
        mem_do_rinst <= !decoder_trigger && !do_waitirq;
        mem_wordsize <= 0;

        current_pc = reg_next_pc;

        (* parallel_case *)
        case (1'b1)
          latched_branch: begin
            current_pc = latched_store ? (latched_stalu ? alu_out_q : reg_out) & ~1 : reg_next_pc;
          end
          latched_store && !latched_branch: begin
          end
          ENABLE_IRQ && irq_state[0]: begin
            current_pc = PROGADDR_IRQ;
            irq_active <= 1;
            mem_do_rinst <= 1;
          end
          ENABLE_IRQ && irq_state[1]: begin
            eoi <= irq_pending & ~irq_mask;
            next_irq_pending = next_irq_pending & irq_mask;
          end
        endcase

        if (ENABLE_TRACE && latched_trace) begin
          latched_trace <= 0;
          trace_valid <= 1;
          if (latched_branch)
            trace_data <= (irq_active ? TRACE_IRQ : 0) | TRACE_BRANCH | (current_pc & 32'hfffffffe);
          else
            trace_data <= (irq_active ? TRACE_IRQ : 0) | (latched_stalu ? alu_out_q : reg_out);
        end

        reg_pc <= current_pc;
        reg_next_pc <= current_pc;

        latched_store <= 0;
        latched_stalu <= 0;
        latched_branch <= 0;
        latched_is_lu <= 0;
        latched_is_lh <= 0;
        latched_is_lb <= 0;
        latched_rd <= decoded_rd;
        // latched_compr <= compressed_instr;

        if (ENABLE_IRQ && ((decoder_trigger && !irq_active && !irq_delay && |(irq_pending & ~irq_mask)) || irq_state)) begin
          irq_state <=
            irq_state == 2'b00 ? 2'b01 :
            irq_state == 2'b01 ? 2'b10 : 2'b00;
          if (ENABLE_IRQ_QREGS)
            latched_rd <= irqregs_offset | irq_state[0];
          else
            latched_rd <= irq_state[0] ? 4 : 3;
        end else
        if (ENABLE_IRQ && (decoder_trigger || do_waitirq) && instr_waitirq) begin
          if (irq_pending) begin
            latched_store <= 1;
            reg_out <= irq_pending;
            reg_next_pc <= current_pc + 4;
            mem_do_rinst <= 1;
          end else
            do_waitirq <= 1;
        end else
        if (decoder_trigger) begin
          irq_delay <= irq_active;
          reg_next_pc <= current_pc + 4;
          if (ENABLE_TRACE)
            latched_trace <= 1;
          if (ENABLE_COUNTERS) begin
            count_instr <= count_instr + 1;
            if (!ENABLE_COUNTERS64) count_instr[63:32] <= 0;
          end
          if (instr_jal) begin
            mem_do_rinst <= 1;
            reg_next_pc <= current_pc + decoded_imm_j;
            latched_branch <= 1;
          end else begin
            mem_do_rinst <= 0;
            mem_do_prefetch <= !instr_jalr && !instr_retirq;
            cpu_state <= cpu_state_ld_rs1;
          end
        end
      end

      cpu_state_ld_rs1: begin
        reg_op1 <= 'bx;
        reg_op2 <= 'bx;

        (* parallel_case *)
        case (1'b1)
          //* error instruction, cause irq_ebreak;
          CATCH_ILLINSN && instr_trap: begin
            if (ENABLE_IRQ && !irq_mask[irq_ebreak] && !irq_active) begin
              next_irq_pending[irq_ebreak] = 1;
              cpu_state <= cpu_state_fetch;
            end else
              cpu_state <= cpu_state_trap;
          end
          ENABLE_COUNTERS && is_rdcycle_rdcycleh_rdinstr_rdinstrh: begin
            (* parallel_case, full_case *)
            case (1'b1)
              instr_rdcycle:
                reg_out <= count_cycle[31:0];
              instr_rdcycleh && ENABLE_COUNTERS64:
                reg_out <= count_cycle[63:32];
              instr_rdinstr:
                reg_out <= count_instr[31:0];
              instr_rdinstrh && ENABLE_COUNTERS64:
                reg_out <= count_instr[63:32];
            endcase
            latched_store <= 1;
            cpu_state <= cpu_state_fetch;
          end
          is_lui_auipc_jal: begin
            reg_op1 <= instr_lui ? 0 : reg_pc;
            reg_op2 <= decoded_imm;
            if (TWO_CYCLE_ALU)
              alu_wait <= 1;
            else
              mem_do_rinst <= mem_do_prefetch;
            cpu_state <= cpu_state_exec;
          end
          ENABLE_IRQ && ENABLE_IRQ_QREGS && instr_getq: begin
            reg_out <= cpuregs_rs1;
            latched_store <= 1;
            cpu_state <= cpu_state_fetch;
          end
          ENABLE_IRQ && ENABLE_IRQ_QREGS && instr_setq: begin
            reg_out <= cpuregs_rs1;
            latched_rd <= latched_rd | irqregs_offset;
            latched_store <= 1;
            cpu_state <= cpu_state_fetch;
          end
          ENABLE_IRQ && instr_retirq: begin
            irq_on <= 1;
            eoi <= 0;
            irq_active <= 0;
            latched_branch <= 1;
            latched_store <= 1;
            reg_out <= CATCH_MISALIGN ? (cpuregs_rs1 & 32'h fffffffe) : cpuregs_rs1;
            cpu_state <= cpu_state_fetch;
          end
          ENABLE_IRQ && instr_maskirq: begin
            latched_store <= 1;
            reg_out <= irq_mask;
            irq_mask <= cpuregs_rs1 | MASKED_IRQ;
            cpu_state <= cpu_state_fetch;
          end
          ENABLE_IRQ && instr_ctlirq: begin
            latched_store <= 1;
            reg_out <= irq_on;
            irq_on <= cpuregs_rs1 & 32'h 0000_0001;
            cpu_state <= cpu_state_fetch;
          end
          ENABLE_IRQ && ENABLE_IRQ_TIMER && instr_timer: begin
            latched_store <= 1;
            reg_out <= timer;
            timer <= cpuregs_rs1;
            timer_conf <= cpuregs_rs1;          
            cpu_state <= cpu_state_fetch;
          end
          is_lb_lh_lw_lbu_lhu && !instr_trap: begin
            reg_op1 <= cpuregs_rs1;
            cpu_state <= cpu_state_ldmem;
            mem_do_rinst <= 1;
          end
          is_slli_srli_srai && !BARREL_SHIFTER: begin
            reg_op1 <= cpuregs_rs1;
            reg_sh <= decoded_rs2;
            cpu_state <= cpu_state_shift;
          end
          is_jalr_addi_slti_sltiu_xori_ori_andi, is_slli_srli_srai && BARREL_SHIFTER: begin
            reg_op1 <= cpuregs_rs1;
            reg_op2 <= is_slli_srli_srai && BARREL_SHIFTER ? decoded_rs2 : decoded_imm;
            if (TWO_CYCLE_ALU)
              alu_wait <= 1;
            else
              mem_do_rinst <= mem_do_prefetch;
            cpu_state <= cpu_state_exec;
          end
          default: begin
            reg_op1 <= cpuregs_rs1;
            if (ENABLE_REGS_DUALPORT) begin
              reg_sh <= cpuregs_rs2;
              reg_op2 <= cpuregs_rs2;
              (* parallel_case *)
              case (1'b1)
                is_sb_sh_sw: begin
                  cpu_state <= cpu_state_stmem;
                  mem_do_rinst <= 1;
                end
                is_sll_srl_sra && !BARREL_SHIFTER: begin
                  cpu_state <= cpu_state_shift;
                end
                default: begin
                  if (TWO_CYCLE_ALU || (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu)) begin
                    alu_wait_2 <= TWO_CYCLE_ALU && (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu);
                    alu_wait <= 1;
                  end else
                    mem_do_rinst <= mem_do_prefetch;
                  cpu_state <= cpu_state_exec;
                end
              endcase
            end else
              cpu_state <= cpu_state_ld_rs2;
          end
        endcase
      end

      cpu_state_ld_rs2: begin
        reg_sh <= cpuregs_rs2;
        reg_op2 <= cpuregs_rs2;

        (* parallel_case *)
        case (1'b1)
          is_sb_sh_sw: begin
            cpu_state <= cpu_state_stmem;
            mem_do_rinst <= 1;
          end
          is_sll_srl_sra && !BARREL_SHIFTER: begin
            cpu_state <= cpu_state_shift;
          end
          default: begin
            if (TWO_CYCLE_ALU || (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu)) begin
              alu_wait_2 <= TWO_CYCLE_ALU && (TWO_CYCLE_COMPARE && is_beq_bne_blt_bge_bltu_bgeu);
              alu_wait <= 1;
            end else
              mem_do_rinst <= mem_do_prefetch;
            cpu_state <= cpu_state_exec;
          end
        endcase
      end

      cpu_state_exec: begin
        reg_out <= reg_pc + decoded_imm;  //* for branch instruction;
        if ((TWO_CYCLE_ALU || TWO_CYCLE_COMPARE) && (alu_wait || alu_wait_2)) begin
          mem_do_rinst <= mem_do_prefetch && !alu_wait_2;
          alu_wait <= alu_wait_2;
        end else
        if (is_beq_bne_blt_bge_bltu_bgeu) begin
          latched_rd <= 0;
          latched_store <= TWO_CYCLE_COMPARE ? alu_out_0_q : alu_out_0;
          latched_branch <= TWO_CYCLE_COMPARE ? alu_out_0_q : alu_out_0;
          if (mem_done)
            cpu_state <= cpu_state_fetch;
          if (TWO_CYCLE_COMPARE ? alu_out_0_q : alu_out_0) begin
            decoder_trigger <= 0;
            set_mem_do_rinst = 1;
          end
        end else begin
          latched_branch <= instr_jalr;
          latched_store <= 1;
          latched_stalu <= 1;
          cpu_state <= cpu_state_fetch;
        end
      end

      cpu_state_shift: begin
        latched_store <= 1;
        if (reg_sh == 0) begin
          reg_out <= reg_op1;
          mem_do_rinst <= mem_do_prefetch;
          cpu_state <= cpu_state_fetch;
        end else if (TWO_STAGE_SHIFT && reg_sh >= 4) begin
          (* parallel_case, full_case *)
          case (1'b1)
            instr_slli || instr_sll: reg_op1 <= reg_op1 << 4;
            instr_srli || instr_srl: reg_op1 <= reg_op1 >> 4;
            instr_srai || instr_sra: reg_op1 <= $signed(reg_op1) >>> 4;
          endcase
          reg_sh <= reg_sh - 4;
        end else begin
          (* parallel_case, full_case *)
          case (1'b1)
            instr_slli || instr_sll: reg_op1 <= reg_op1 << 1;
            instr_srli || instr_srl: reg_op1 <= reg_op1 >> 1;
            instr_srai || instr_sra: reg_op1 <= $signed(reg_op1) >>> 1;
          endcase
          reg_sh <= reg_sh - 1;
        end
      end

      cpu_state_stmem: begin
        if (ENABLE_TRACE)
          reg_out <= reg_op2;
        if (!mem_do_prefetch || mem_done) begin
          if (!mem_do_wdata) begin
            (* parallel_case, full_case *)
            case (1'b1)
              instr_sb: mem_wordsize <= 2;
              instr_sh: mem_wordsize <= 1;
              instr_sw: mem_wordsize <= 0;
            endcase
            if (ENABLE_TRACE) begin
              trace_valid <= 1;
              trace_data <= (irq_active ? TRACE_IRQ : 0) | TRACE_ADDR | ((reg_op1 + decoded_imm) & 32'hffffffff);
            end
            reg_op1 <= reg_op1 + decoded_imm;
            set_mem_do_wdata = 1;
          end
          if (!mem_do_prefetch && mem_done) begin
            cpu_state <= cpu_state_fetch;
            decoder_trigger <= 1;
            decoder_pseudo_trigger <= 1;
          end
        end
      end

      cpu_state_ldmem: begin
        latched_store <= 1;
        if (!mem_do_prefetch || mem_done) begin
          if (!mem_do_rdata) begin
            (* parallel_case, full_case *)
            case (1'b1)
              instr_lb || instr_lbu: mem_wordsize <= 2;
              instr_lh || instr_lhu: mem_wordsize <= 1;
              instr_lw: mem_wordsize <= 0;
            endcase
            latched_is_lu <= is_lbu_lhu_lw;
            latched_is_lh <= instr_lh;
            latched_is_lb <= instr_lb;
            if (ENABLE_TRACE) begin
              trace_valid <= 1;
              trace_data <= (irq_active ? TRACE_IRQ : 0) | TRACE_ADDR | ((reg_op1 + decoded_imm) & 32'hffffffff);
            end
            reg_op1 <= reg_op1 + decoded_imm;
            set_mem_do_rdata = 1;
          end
          if (!mem_do_prefetch && mem_done) begin
            (* parallel_case, full_case *)
            case (1'b1)
              latched_is_lu: reg_out <= mem_rdata_word;
              latched_is_lh: reg_out <= $signed(mem_rdata_word[15:0]);
              latched_is_lb: reg_out <= $signed(mem_rdata_word[7:0]);
            endcase
            decoder_trigger <= 1;
            decoder_pseudo_trigger <= 1;
            cpu_state <= cpu_state_fetch;
          end
        end
      end
    endcase

    if (CATCH_MISALIGN && resetn && (mem_do_rdata || mem_do_wdata)) begin
      if (mem_wordsize == 0 && reg_op1[1:0] != 0) begin
        if (ENABLE_IRQ && !irq_mask[irq_buserror] && !irq_active) begin
          next_irq_pending[irq_buserror] = 1;
        end else
          cpu_state <= cpu_state_trap;
      end
      if (mem_wordsize == 1 && reg_op1[0] != 0) begin
        if (ENABLE_IRQ && !irq_mask[irq_buserror] && !irq_active) begin
          next_irq_pending[irq_buserror] = 1;
        end else
          cpu_state <= cpu_state_trap;
      end
    end
    if (CATCH_MISALIGN && resetn && mem_do_rinst && (|reg_pc[1:0])) begin
      if (ENABLE_IRQ && !irq_mask[irq_buserror] && !irq_active) begin
        next_irq_pending[irq_buserror] = 1;
      end else
        cpu_state <= cpu_state_trap;
    end
    if (!CATCH_ILLINSN && decoder_trigger_q && !decoder_pseudo_trigger_q && instr_ecall_ebreak) begin
      cpu_state <= cpu_state_trap;
    end

    if (!resetn || mem_done) begin
      mem_do_prefetch <= 0;
      mem_do_rinst <= 0;
      mem_do_rdata <= 0;
      mem_do_wdata <= 0;
    end

    if (set_mem_do_rinst)
      mem_do_rinst <= 1;
    if (set_mem_do_rdata)
      mem_do_rdata <= 1;
    if (set_mem_do_wdata)
      mem_do_wdata <= 1;

    irq_pending <= irq_on ? next_irq_pending & ~MASKED_IRQ: next_irq_pending & ~SYS_MASKED_IRQ;

    if (!CATCH_MISALIGN) begin
      reg_pc[1:0] <= 0;
      reg_next_pc[1:0] <= 0;
    end
    current_pc = 'bx;
  end


  // Formal Verification

endmodule
