 /*
 *  picoSoC_hardware -- SoC Hardware for RISCV-32I core.
 *
 *  Copyright (C) 2021-2022 Junnan Li <lijunnan@nudt.edu.cn>.
 *  Copyright and related rights are licensed under the MIT license.
 *
 *  Date: 2022.02.20
 *  Description: This module is used to process packets by CPU.
 */

`timescale 1 ns / 1 ps

module memPkt(
  input               clk,
  input               rst_n,

  input               data_in_valid,  // input data valid
  input       [133:0] data_in,    

  output  reg         data_out_valid, // output data valid
  (* mark_debug = "true"*)output  reg [133:0] data_out,       // output data

  input               memPkt_rden,    // mem interface
  input               memPkt_wren,
  input       [31:0]  memPkt_addr,
  input       [31:0]  memPkt_wdata,
  input       [3:0]   memPkt_wstrb,
  output  reg [31:0]  memPkt_rdata,
  output  reg         memPkt_ready 
);


/** state_sendPkt is used to out pkt generated by CPU;
 */
reg       state_sendPkt;
parameter IDLE_S      = 1'd0,
          WAIT_TAIL_S = 1'd1;

/** fifo signals;
 */
(* mark_debug = "true"*)reg   [133:0] din_pktRecv, din_pktSend;
(* mark_debug = "true"*)reg           wren_pktRecv, wren_pktSend;
(* mark_debug = "true"*)reg           rden_pktRecv, rden_pktSend;
(* mark_debug = "true"*)wire  [133:0] dout_pktRecv, dout_pktSend;
(* mark_debug = "true"*)wire          empty_pktRecv, empty_pktSend;

/** cnt_rden_last8b/cnt_wren_last8b is used to count times that C program has
 *    read/written the last 8b data, to change 128b recvPkt_reg/sendPkt_reg;
 *  recvPkt_reg/sendPkt_reg is 128b, used for C program to read/write;
 *  length is 16b, record pkt's length (in B);
 *  tag is 2b, "tag[0]=1" -> recv pkt (finish); "tag[0]=2" -> finish read;
 *             "tag[1]=1" -> finish writing; "tag[1]=2" -> send pkt (finish);
 *    tag[0] is operated by hw, while tag[1] is operated by CUP;
 *  temp_sendTag used to delay sending pkt, we meet mistake when sending just 
 *    after writing tag;
 */
(* mark_debug = "true"*)reg   [1:0]   cnt_rden_last8b, cnt_wren_last8b;
(* mark_debug = "true"*)reg   [127:0] recvPkt_reg, sendPkt_reg;
(* mark_debug = "true"*)reg   [15:0]  length[1:0];  //* 0 is recv, 1 is send;
(* mark_debug = "true"*)reg   [7:0]   sendLength;
(* mark_debug = "true"*)reg   [1:0]   tag[1:0];     //* 0 is recv, 1 is send;
(* mark_debug = "true"*)reg   [3:0]   temp_sendTag; //* meet mistake when sending just after writing tag;

/** state machine for write recv pkt from fifo to reg, or write sending 
*   pkt from reg to fifo;
*     1) fifo just buffer one pkt;
*     2) read one pkt data after reading the last 8b;
*     3) write one pkt data after writing the last 8b;
*/
always @(posedge clk or negedge rst_n) begin
  if (!rst_n) begin
    // reset
    memPkt_rdata          <= 32'b0;   //* mem interface (output);
    memPkt_ready          <= 1'b0;
    din_pktRecv           <= 134'b0;  //* fifo interface;
    wren_pktRecv          <= 1'b0;
    din_pktSend           <= {2'b10,132'b0};
    wren_pktSend          <= 1'b0;
    rden_pktRecv          <= 1'b0;
    rden_pktSend          <= 1'b0;   
    cnt_rden_last8b       <= 2'd0;    //* count info;
    cnt_wren_last8b       <= 2'd0;
    recvPkt_reg           <= 128'b0;  //* reg to read/write;
    sendPkt_reg           <= 128'b0;
    {length[1],length[0]} <= 32'b0;
    sendLength            <= 8'b0;
    {tag[1],tag[0]}       <= 4'b0;
    temp_sendTag          <= 4'b0;    //* delay sending;

    data_out_valid        <= 1'b0;    //* pkt out;
    data_out              <= 134'b0;
    state_sendPkt         <= IDLE_S;
  end
  else begin
    //* 1) recv pkt (write fifo_recv), and calculate length;
    //* 2) discard CPU configuration packets (0x90..);
      din_pktRecv           <= data_in;
      if(data_in_valid == 1'b1 && data_in[133:132] == 2'b01 &&
        data_in[31:24] != 8'h90 && tag[0][0] == 1'b0) 
      begin
        wren_pktRecv        <= 1'b1;
        length[0]           <= 16'b0;
      end
      else begin
        wren_pktRecv        <= wren_pktRecv & data_in_valid;
        length[0]           <= (wren_pktRecv == 1'b1)? (length[0] + 16'd1 + 
                                  {12'b0, din_pktRecv[131:128]}): length[0];
      end

    //* write recv pkt from fifo to reg, big-end <-> small-end:
    //*   1) C program has finished reading current packet, i.e., tag[0][0] == 1'b0;
    //*   2) C program has finished reading current 128b data; 
      rden_pktRecv          <= 1'b0;
      if((tag[0][0] == 1'b0 && empty_pktRecv == 1'b0 && wren_pktRecv == 1'b0)) begin 
        tag[0][0]           <= 1'd1;
        rden_pktRecv        <= 1'b1;
        recvPkt_reg         <= {dout_pktRecv[96+:8],dout_pktRecv[104+:8],
                                dout_pktRecv[112+:8],dout_pktRecv[120+:8],
                                dout_pktRecv[64+:8],dout_pktRecv[72+:8],
                                dout_pktRecv[80+:8],dout_pktRecv[88+:8],
                                dout_pktRecv[32+:8],dout_pktRecv[40+:8],
                                dout_pktRecv[48+:8],dout_pktRecv[56+:8],
                                dout_pktRecv[0+:8],dout_pktRecv[8+:8],
                                dout_pktRecv[16+:8],dout_pktRecv[24+:8]};
      end
      else if(memPkt_rden == 1'b1 && cnt_rden_last8b == 2'd3 && 
        memPkt_addr[31:24] == 8'h12 && empty_pktRecv == 1'b0) 
      begin
        rden_pktRecv        <= 1'b1;
        recvPkt_reg         <= {dout_pktRecv[96+:8],dout_pktRecv[104+:8],
                                dout_pktRecv[112+:8],dout_pktRecv[120+:8],
                                dout_pktRecv[64+:8],dout_pktRecv[72+:8],
                                dout_pktRecv[80+:8],dout_pktRecv[88+:8],
                                dout_pktRecv[32+:8],dout_pktRecv[40+:8],
                                dout_pktRecv[48+:8],dout_pktRecv[56+:8],
                                dout_pktRecv[0+:8],dout_pktRecv[8+:8],
                                dout_pktRecv[16+:8],dout_pktRecv[24+:8]};
      end
      else if(tag[0][1] == 1'b1) begin //* clear tag[0][0], e.g., recv pkt isn't ready;
        tag[0][0]           <= 1'd0;
      end
    
    //* update cnt_rden_last8b;
      if(memPkt_rden == 1'b1 && memPkt_addr[31:24] == 8'h12) begin
        cnt_rden_last8b     <= (memPkt_addr[3:2] == 2'h1)? (cnt_rden_last8b + 2'd1): 2'd0;
      end

    //* 1) send pkt, i.e., C program has finished writing packet (tag[1][0] == 1'd1);
    //* 2) delay 4 clock sending, since meet mistake when sending just after writing tag;
      temp_sendTag          <= {temp_sendTag[2:0],tag[1][0]};
      case(state_sendPkt)
        IDLE_S: begin
          data_out_valid    <= 1'b0;
          if(temp_sendTag[3] == 1'd1 && empty_pktSend == 1'b0) begin
            rden_pktSend    <= 1'b1;
            state_sendPkt   <= WAIT_TAIL_S;
          end
        end
        WAIT_TAIL_S: begin
          data_out_valid    <= 1'b1;
          data_out          <= dout_pktSend;
          if(dout_pktSend[133:132] == 2'b10) begin
            rden_pktSend    <= 1'b0;
            state_sendPkt   <= IDLE_S;
          end
        end
        default: begin
          state_sendPkt     <= IDLE_S;
        end
      endcase
    
    //* write send pkt from reg to fifo, big-end <-> small-end:
    //*   1) C program has finished writing current packet, i.e., tag[1] == 2'b1;
    //*   2) C program has finished writing current 128b data, but not last 128b data;
      wren_pktSend          <= 1'b0;
      if(tag[1] == 2'd1) begin //* one pkt is ready;
        wren_pktSend        <= 1'b1;
        din_pktSend[127:0]  <= {sendPkt_reg[96+:8], sendPkt_reg[104+:8],
                                sendPkt_reg[112+:8],sendPkt_reg[120+:8],
                                sendPkt_reg[64+:8], sendPkt_reg[72+:8],
                                sendPkt_reg[80+:8], sendPkt_reg[88+:8],
                                sendPkt_reg[32+:8], sendPkt_reg[40+:8],
                                sendPkt_reg[48+:8], sendPkt_reg[56+:8],
                                sendPkt_reg[0+:8],  sendPkt_reg[8+:8],
                                sendPkt_reg[16+:8], sendPkt_reg[24+:8]};
        din_pktSend[133:132]  <= 2'b10;
        din_pktSend[131:128]  <= length[1][3:0] - 4'd1;
      end
      else if(memPkt_wren == 1'b1 && cnt_wren_last8b == 2'd3 && 
        memPkt_addr[31:24] == 8'h11 && memPkt_addr[3:2] == 2'h1) 
      begin
        sendLength          <= sendLength - 8'd1;
        wren_pktSend        <= (|{sendLength,length[1][3:0]})? 1'b1:1'b0;
        din_pktSend[127:0]  <= {sendPkt_reg[96+:8], sendPkt_reg[104+:8],
                                sendPkt_reg[112+:8],sendPkt_reg[120+:8],
                                sendPkt_reg[64+:8], sendPkt_reg[72+:8],
                                sendPkt_reg[80+:8], sendPkt_reg[88+:8],
                                sendPkt_reg[32+:8], sendPkt_reg[40+:8],
                                sendPkt_reg[48+:8], sendPkt_reg[56+:8],
                                sendPkt_reg[0+:8],  sendPkt_reg[8+:8],
                                sendPkt_reg[16+:8], memPkt_wdata[7:0]};
        din_pktSend[133:132]  <= (din_pktSend[133:132] == 2'b10)? 2'd1: 2'd0;
        din_pktSend[131:128]  <= 4'hf;
      end
      else if(memPkt_wren == 1'b1 && memPkt_addr[10:2] == 9'd1 && 
        memPkt_addr[31:24] == 8'h11) 
      begin
        sendLength          <= memPkt_wdata[11:4] - 8'd1;
      end
    
    //* update cnt_rden_last8b;
      if(memPkt_wren == 1'b1 && memPkt_addr[31:24] == 8'h11) begin
        cnt_wren_last8b     <= (memPkt_addr[3:2] == 2'h1)? (cnt_wren_last8b + 2'd1): 2'd0;
      end
    
    //* proc pkt;
    //*   1) read pkt data;
      tag[1]                <= 2'b0;
      tag[0][1]             <= 1'b0;
      sendPkt_reg           <= sendPkt_reg;
      if(memPkt_rden == 1'b1 && memPkt_addr[31:24] == 8'h12) begin
        memPkt_ready        <= 1'b1;
        if(memPkt_addr[10:3] == 8'b0)
          memPkt_rdata      <= (memPkt_addr[2] == 1'b0)? {30'b0,tag[0]}: {16'b0,length[0]};
        else begin
          (*full_case, parallel_case*)
          case(memPkt_addr[3:2])
            2'd0: memPkt_rdata  <= recvPkt_reg[32+:32];
            2'd1: memPkt_rdata  <= recvPkt_reg[0+:32];
            2'd2: memPkt_rdata  <= recvPkt_reg[96+:32];
            2'd3: memPkt_rdata  <= recvPkt_reg[64+:32];
          endcase
        end
      end
    //*   2) write pkt data;
      else if(memPkt_wren == 1'b1 && memPkt_addr[31:24] == 8'h11) begin
        memPkt_ready        <= 1'b1;
        if(memPkt_addr[10:3] == 8'b0) begin
          tag[1]            <= (memPkt_addr[2] == 1'b0)? memPkt_wdata[1:0]:  tag[1];
          length[1]         <= (memPkt_addr[2] == 1'b1)? memPkt_wdata[15:0]: length[1];
        end
        else begin
          (*full_case, parallel_case*)
          case(memPkt_addr[3:2])
            2'd0: begin
              if (memPkt_wstrb[0]) sendPkt_reg[32*1+7:32*1]     <= memPkt_wdata[ 7: 0];
              if (memPkt_wstrb[1]) sendPkt_reg[32*1+15:32*1+8]  <= memPkt_wdata[15: 8];
              if (memPkt_wstrb[2]) sendPkt_reg[32*1+23:32*1+16] <= memPkt_wdata[23:16];
              if (memPkt_wstrb[3]) sendPkt_reg[32*1+31:32*1+24] <= memPkt_wdata[31:24];
            end
            2'd1: begin
              if (memPkt_wstrb[0]) sendPkt_reg[32*0+7:32*0]     <= memPkt_wdata[ 7: 0];
              if (memPkt_wstrb[1]) sendPkt_reg[32*0+15:32*0+8]  <= memPkt_wdata[15: 8];
              if (memPkt_wstrb[2]) sendPkt_reg[32*0+23:32*0+16] <= memPkt_wdata[23:16];
              if (memPkt_wstrb[3]) sendPkt_reg[32*0+31:32*0+24] <= memPkt_wdata[31:24];
            end
            2'd2: begin
              if (memPkt_wstrb[0]) sendPkt_reg[32*3+7:32*3]     <= memPkt_wdata[ 7: 0];
              if (memPkt_wstrb[1]) sendPkt_reg[32*3+15:32*3+8]  <= memPkt_wdata[15: 8];
              if (memPkt_wstrb[2]) sendPkt_reg[32*3+23:32*3+16] <= memPkt_wdata[23:16];
              if (memPkt_wstrb[3]) sendPkt_reg[32*3+31:32*3+24] <= memPkt_wdata[31:24];
            end
            2'd3: begin
              if (memPkt_wstrb[0]) sendPkt_reg[32*2+7:32*2]     <= memPkt_wdata[ 7: 0];
              if (memPkt_wstrb[1]) sendPkt_reg[32*2+15:32*2+8]  <= memPkt_wdata[15: 8];
              if (memPkt_wstrb[2]) sendPkt_reg[32*2+23:32*2+16] <= memPkt_wdata[23:16];
              if (memPkt_wstrb[3]) sendPkt_reg[32*2+31:32*2+24] <= memPkt_wdata[31:24];
            end
          endcase
        end
      end
    //*   3) read tag[1], or other address (return 0);
      else if(memPkt_rden == 1'b1 && memPkt_addr[31:24] == 8'h11) begin
        memPkt_ready        <= 1'b1;
        if(memPkt_addr[10:2] == 9'b0) memPkt_rdata  <= 32'd2;
        else                          memPkt_rdata  <= 32'd0;
      end
    //*   4) write tag[0], or other address (nop);
      else if(memPkt_wren == 1'b1 && memPkt_addr[31:24] == 8'h12) begin
        memPkt_ready        <= 1'b1;
        if(memPkt_addr[10:2] == 9'b0) tag[0][1]     <= 1'd1;
      end
      else
        memPkt_ready        <= 1'b0;
  end
end




/** fifo used to buffer recv/send pkt*/
fifo_134b_512 fifo_pktRecv (
  .clk(clk),              // input wire clk
  .srst(!rst_n),          // input wire srst
  .din(din_pktRecv),      // input wire [133 : 0] din
  .wr_en(wren_pktRecv),   // input wire wr_en
  .rd_en(rden_pktRecv),   // input wire rd_en
  .dout(dout_pktRecv),    // output wire [133 : 0] dout
  .full(),                // output wire full
  .empty(empty_pktRecv)   // output wire empty
);

fifo_134b_512 fifo_pktSend (
  .clk(clk),              // input wire clk
  .srst(!rst_n),          // input wire srst
  .din(din_pktSend),      // input wire [133 : 0] din
  .wr_en(wren_pktSend),   // input wire wr_en
  .rd_en(rden_pktSend),   // input wire rd_en
  .dout(dout_pktSend),    // output wire [133 : 0] dout
  .full(),                // output wire full
  .empty(empty_pktSend)   // output wire empty
);




endmodule
